<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-64.0627,6.74441,310.561,-188.574</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>101,-18.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>87,-19</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_INVERTER</type>
<position>93.5,-23</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_INVERTER</type>
<position>107.5,-22.5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_AND2</type>
<position>118.5,-32.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>103,-13.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>86.5,-13</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>66,-13.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>51.5,-13.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>35,-13.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>23,-13.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>1.5,-13.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>-14,-13.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND2</type>
<position>118.5,-41</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>65.5,-18.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>51.5,-18.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_INVERTER</type>
<position>55.5,-23</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_INVERTER</type>
<position>69.5,-23</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>118.5,-55.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>118.5,-64</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>36.5,-18.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>22.5,-18.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_INVERTER</type>
<position>26.5,-23</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_INVERTER</type>
<position>40.5,-23</position>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND2</type>
<position>119,-77.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND2</type>
<position>119,-85</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>0.5,-19</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>-13.5,-19</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_INVERTER</type>
<position>-9.5,-23.5</position>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_INVERTER</type>
<position>4.5,-23.5</position>
<input>
<ID>IN_0</ID>25 </input>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>119,-100.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_AND2</type>
<position>119,-108.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_OR4</type>
<position>200,-55.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>53 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>61 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_OR4</type>
<position>199.5,-81</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>62 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND4</type>
<position>199.5,-141</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>51 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>227,-141.5</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>BE_NOR2</type>
<position>128.5,-36.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>BE_NOR2</type>
<position>129.5,-59.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>BE_NOR2</type>
<position>130,-81.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>BE_NOR2</type>
<position>130,-104.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>161,-50.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_AND2</type>
<position>161,-63</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_AND3</type>
<position>160.5,-72.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>45 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>217,-81</position>
<input>
<ID>N_in0</ID>57 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>GA_LED</type>
<position>212,-55.5</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_AND3</type>
<position>160.5,-86.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>46 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_AND4</type>
<position>160.5,-99</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>51 </input>
<input>
<ID>IN_3</ID>47 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND4</type>
<position>160,-118.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>51 </input>
<input>
<ID>IN_3</ID>48 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-33.5,87,-21</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-33.5 1</intersection>
<intersection>-23 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-33.5,115.5,-33.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>87,-23,90.5,-23</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-42,101,-20.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-42 3</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101,-22.5,104.5,-22.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>101 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101,-42,115.5,-42</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-31.5,113,-22.5</points>
<intersection>-31.5 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,-31.5,115.5,-31.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>113 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-22.5,113,-22.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>113 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-40,98,-23</points>
<intersection>-40 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-40,115.5,-40</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-23,98,-23</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-56.5,51.5,-20.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>-56.5 1</intersection>
<intersection>-23 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-56.5,115.5,-56.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>51.5,-23,52.5,-23</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-65,65.5,-20.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>-65 3</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-23,66.5,-23</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>65.5,-65,115.5,-65</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-54.5,74,-23</points>
<intersection>-54.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-54.5,115.5,-54.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-23,74,-23</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-63,115.5,-63</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>58.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58.5,-63,58.5,-23</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-63 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-78.5,22.5,-20.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 1</intersection>
<intersection>-23 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-78.5,116,-78.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>22.5,-23,23.5,-23</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-86,36.5,-20.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>-86 3</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-23,37.5,-23</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36.5,-86,116,-86</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-76.5,45,-23</points>
<intersection>-76.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-76.5,116,-76.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-23,45,-23</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-84,116,-84</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>29.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29.5,-84,29.5,-23</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>-84 1</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-101.5,-13.5,-21</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-101.5 1</intersection>
<intersection>-23.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-101.5,116,-101.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-13.5,-23.5,-12.5,-23.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-109.5,0.5,-21</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-109.5 3</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-23.5,1.5,-23.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>0.5,-109.5,116,-109.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-99.5,9,-23.5</points>
<intersection>-99.5 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-99.5,116,-99.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-23.5,9,-23.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-107.5,116,-107.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-6.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-6.5,-107.5,-6.5,-23.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>-107.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>202.5,-141,226,-141</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>226 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>226,-141.5,226,-141</points>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<intersection>-141 1</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-35.5,125.5,-27.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-35.5 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-27.5,197,-27.5</points>
<intersection>125.5 0</intersection>
<intersection>197 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-35.5,125.5,-35.5</points>
<intersection>121.5 4</intersection>
<intersection>125.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>197,-52.5,197,-27.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>121.5,-35.5,121.5,-32.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>-35.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-44,125,-37.5</points>
<intersection>-44 3</intersection>
<intersection>-41 1</intersection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-41,125,-41</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-37.5,125.5,-37.5</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>125,-44,152.5,-44</points>
<intersection>125 0</intersection>
<intersection>152.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>152.5,-80,152.5,-44</points>
<intersection>-80 5</intersection>
<intersection>-44 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>152.5,-80,196.5,-80</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>152.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-58.5,124,-51.5</points>
<intersection>-58.5 5</intersection>
<intersection>-55.5 1</intersection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-55.5,124,-55.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124,-51.5,158,-51.5</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>124,-58.5,126.5,-58.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-64,124,-60.5</points>
<intersection>-64 1</intersection>
<intersection>-60.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-64,158,-64</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>124,-60.5,126.5,-60.5</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>124 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-80.5,124.5,-74.5</points>
<intersection>-80.5 3</intersection>
<intersection>-77.5 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-77.5,124.5,-77.5</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-74.5,157.5,-74.5</points>
<connection>
<GID>85</GID>
<name>IN_2</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>124.5,-80.5,127,-80.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-88.5,125,-82.5</points>
<intersection>-88.5 2</intersection>
<intersection>-85 1</intersection>
<intersection>-82.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-85,125,-85</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-88.5,157.5,-88.5</points>
<connection>
<GID>88</GID>
<name>IN_2</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>125,-82.5,127,-82.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-102,124.5,-100.5</points>
<intersection>-102 2</intersection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-100.5,124.5,-100.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-102,157.5,-102</points>
<connection>
<GID>90</GID>
<name>IN_3</name></connection>
<intersection>124.5 0</intersection>
<intersection>127 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127,-103.5,127,-102</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-102 2</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-108.5,124.5,-105.5</points>
<intersection>-108.5 1</intersection>
<intersection>-105.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-108.5,124.5,-108.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-105.5,127,-105.5</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>124.5 0</intersection>
<intersection>127 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>127,-121.5,127,-105.5</points>
<intersection>-121.5 4</intersection>
<intersection>-105.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>127,-121.5,157,-121.5</points>
<connection>
<GID>91</GID>
<name>IN_3</name></connection>
<intersection>127 3</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-138,150.5,-36.5</points>
<intersection>-138 1</intersection>
<intersection>-115.5 8</intersection>
<intersection>-96 7</intersection>
<intersection>-84.5 6</intersection>
<intersection>-70.5 5</intersection>
<intersection>-62 4</intersection>
<intersection>-49.5 3</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-138,196.5,-138</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131.5,-36.5,150.5,-36.5</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>150.5,-49.5,158,-49.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>150.5,-62,158,-62</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>150.5,-70.5,157.5,-70.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>150.5,-84.5,157.5,-84.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>150.5,-96,157.5,-96</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>150.5,-115.5,157,-115.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>150.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-140,148.5,-59.5</points>
<intersection>-140 1</intersection>
<intersection>-117.5 6</intersection>
<intersection>-98 5</intersection>
<intersection>-86.5 4</intersection>
<intersection>-72.5 3</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148.5,-140,196.5,-140</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-59.5,148.5,-59.5</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148.5,-72.5,157.5,-72.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>148.5,-86.5,157.5,-86.5</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>148.5,-98,157.5,-98</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>148.5,-117.5,157,-117.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147,-142,147,-81.5</points>
<intersection>-142 1</intersection>
<intersection>-119.5 4</intersection>
<intersection>-100 3</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147,-142,196.5,-142</points>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133,-81.5,147,-81.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>147,-100,157.5,-100</points>
<connection>
<GID>90</GID>
<name>IN_2</name></connection>
<intersection>147 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>147,-119.5,157,-119.5</points>
<connection>
<GID>91</GID>
<name>IN_2</name></connection>
<intersection>147 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-144,145.5,-104.5</points>
<intersection>-144 1</intersection>
<intersection>-104.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,-144,196.5,-144</points>
<connection>
<GID>73</GID>
<name>IN_3</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133,-104.5,145.5,-104.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-54.5,179.5,-50.5</points>
<intersection>-54.5 1</intersection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179.5,-54.5,197,-54.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>179.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>164,-50.5,179.5,-50.5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>179.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-78,168,-63</points>
<intersection>-78 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>164,-63,168,-63</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168,-78,196.5,-78</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-55.5,211,-55.5</points>
<connection>
<GID>87</GID>
<name>N_in0</name></connection>
<connection>
<GID>69</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>203.5,-81,216,-81</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,-72.5,180,-56.5</points>
<intersection>-72.5 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180,-56.5,197,-56.5</points>
<connection>
<GID>69</GID>
<name>IN_2</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-72.5,180,-72.5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>180 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-86.5,168,-82</points>
<intersection>-86.5 2</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-82,196.5,-82</points>
<connection>
<GID>71</GID>
<name>IN_2</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-86.5,168,-86.5</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,-99,181,-58.5</points>
<intersection>-99 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181,-58.5,197,-58.5</points>
<connection>
<GID>69</GID>
<name>IN_3</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-99,181,-99</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<intersection>181 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-118.5,183,-84</points>
<intersection>-118.5 2</intersection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-84,196.5,-84</points>
<connection>
<GID>71</GID>
<name>IN_3</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-118.5,183,-118.5</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-140.746,70.741,280.706,-148.992</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>21,27</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>-54.5,30.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_INVERTER</type>
<position>-50.5,26.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_INVERTER</type>
<position>27.5,23</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_AND2</type>
<position>82.5,7</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>21,33</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>-54,36</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>32.5,33</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>-43.5,36</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>42,33</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>-32.5,36</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>54,33</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>-20,36.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>82.5,-1.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>33,27.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>-43.5,31</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_INVERTER</type>
<position>-39.5,26.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_INVERTER</type>
<position>37,23</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_AND2</type>
<position>82.5,-16</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>82.5,-24.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>42,27.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>-33,31</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_INVERTER</type>
<position>-29,26.5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_INVERTER</type>
<position>46,23</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_AND2</type>
<position>83,-38</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>83,-45.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>53,28</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-19.5,31</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_INVERTER</type>
<position>-15.5,26.5</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_INVERTER</type>
<position>57,23</position>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_AND2</type>
<position>83,-61</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND2</type>
<position>83,-69</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_OR4</type>
<position>164,-17</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>67 </input>
<input>
<ID>IN_2</ID>71 </input>
<input>
<ID>IN_3</ID>73 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_OR4</type>
<position>163.5,-41.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>72 </input>
<input>
<ID>IN_3</ID>74 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND4</type>
<position>168.5,-91.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>66 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>68</ID>
<type>GA_LED</type>
<position>185.5,-69.5</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>BE_NOR2</type>
<position>92.5,3</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>BE_NOR2</type>
<position>93.5,-20</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>BE_NOR2</type>
<position>94,-42</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>BE_NOR2</type>
<position>94,-65</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_AND2</type>
<position>125,-11</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_AND2</type>
<position>125,-23.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_AND3</type>
<position>124.5,-33</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>38 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>92</ID>
<type>GA_LED</type>
<position>185.5,-41.5</position>
<input>
<ID>N_in0</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>GA_LED</type>
<position>185.5,-17</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_AND3</type>
<position>124.5,-47</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>39 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_AND4</type>
<position>124.5,-59.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>55 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND4</type>
<position>124,-79</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<input>
<ID>IN_2</ID>65 </input>
<input>
<ID>IN_3</ID>60 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>185.5,-12.5</position>
<gparam>LABEL_TEXT A  B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>186,-64</position>
<gparam>LABEL_TEXT A = B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>186.5,-36.5</position>
<gparam>LABEL_TEXT A > B</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>72.5,29</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>2 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>103</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-1,29.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>5 </input>
<input>
<ID>IN_3</ID>1 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,6,-54.5,28.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>6 1</intersection>
<intersection>12 6</intersection>
<intersection>26.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54.5,6,79.5,6</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-54.5,26.5,-53.5,26.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-54.5,12,-9,12</points>
<intersection>-54.5 0</intersection>
<intersection>-9 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-9,12,-9,31.5</points>
<intersection>12 6</intersection>
<intersection>31.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-9,31.5,-4,31.5</points>
<connection>
<GID>103</GID>
<name>IN_3</name></connection>
<intersection>-9 7</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-2.5,21,25</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-2.5 3</intersection>
<intersection>12.5 7</intersection>
<intersection>23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,23,24.5,23</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>21,-2.5,79.5,-2.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21,12.5,65.5,12.5</points>
<intersection>21 0</intersection>
<intersection>65.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>65.5,12.5,65.5,31</points>
<intersection>12.5 7</intersection>
<intersection>31 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>65.5,31,69.5,31</points>
<connection>
<GID>102</GID>
<name>IN_3</name></connection>
<intersection>65.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,8,79.5,8</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>30.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30.5,8,30.5,23</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>8 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,-0.5,79.5,-0.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-46 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-46,-0.5,-46,26.5</points>
<intersection>-0.5 1</intersection>
<intersection>26.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-47.5,26.5,-46,26.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-46 5</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43.5,-17,-43.5,29</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>-17 1</intersection>
<intersection>14 4</intersection>
<intersection>26.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-43.5,-17,79.5,-17</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-43.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-43.5,14,-7.5,14</points>
<intersection>-43.5 0</intersection>
<intersection>-7.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-7.5,14,-7.5,30.5</points>
<intersection>14 4</intersection>
<intersection>30.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-7.5,30.5,-4,30.5</points>
<connection>
<GID>103</GID>
<name>IN_2</name></connection>
<intersection>-7.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-43.5,26.5,-42.5,26.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-25.5,33,25.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 3</intersection>
<intersection>14 1</intersection>
<intersection>23 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,14,66.5,14</points>
<intersection>33 0</intersection>
<intersection>66.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-25.5,79.5,-25.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>66.5,14,66.5,30</points>
<intersection>14 1</intersection>
<intersection>30 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>33,23,34,23</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>66.5,30,69.5,30</points>
<connection>
<GID>102</GID>
<name>IN_2</name></connection>
<intersection>66.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-15,79.5,-15</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>40 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40,-15,40,23</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-15 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-35.5,-23.5,79.5,-23.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-35.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-35.5,-23.5,-35.5,26.5</points>
<intersection>-23.5 1</intersection>
<intersection>26.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-36.5,26.5,-35.5,26.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-39,-33,29</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-39 1</intersection>
<intersection>17 4</intersection>
<intersection>26.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33,-39,80,-39</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-33 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-33,17,-6.5,17</points>
<intersection>-33 0</intersection>
<intersection>-6.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-6.5,17,-6.5,29.5</points>
<intersection>17 4</intersection>
<intersection>29.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-6.5,29.5,-4,29.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>-6.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-33,26.5,-32,26.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-33 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-46.5,42,25.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>-46.5 3</intersection>
<intersection>15 1</intersection>
<intersection>23 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,15,67.5,15</points>
<intersection>42 0</intersection>
<intersection>67.5 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>42,-46.5,80,-46.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>42 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>67.5,15,67.5,29</points>
<intersection>15 1</intersection>
<intersection>29 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>67.5,29,69.5,29</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>67.5 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>42,23,43,23</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-37,80,-37</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-37,50,23</points>
<intersection>-37 1</intersection>
<intersection>23 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>49,23,50,23</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>50 3</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-24,-44.5,80,-44.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-24 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-24,-44.5,-24,26.5</points>
<intersection>-44.5 1</intersection>
<intersection>26.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-26,26.5,-24,26.5</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-24 8</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-62,-19.5,29</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-62 1</intersection>
<intersection>19.5 4</intersection>
<intersection>26.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19.5,-62,80,-62</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-19.5,19.5,-5,19.5</points>
<intersection>-19.5 0</intersection>
<intersection>-5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-5,19.5,-5,28.5</points>
<intersection>19.5 4</intersection>
<intersection>28.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-19.5,26.5,-18.5,26.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-5,28.5,-4,28.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-5 5</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-70,53,26</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-70 3</intersection>
<intersection>18 1</intersection>
<intersection>23 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,18,68.5,18</points>
<intersection>53 0</intersection>
<intersection>68.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>53,-70,80,-70</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>68.5,18,68.5,28</points>
<intersection>18 1</intersection>
<intersection>28 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>53,23,54,23</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>68.5,28,69.5,28</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>68.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-60,62,23</points>
<intersection>-60 1</intersection>
<intersection>23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-60,80,-60</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,23,62,23</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11,-68,80,-68</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-11 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-11,-68,-11,26.5</points>
<intersection>-68 1</intersection>
<intersection>26.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-12.5,26.5,-11,26.5</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-11 6</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>171.5,-91.5,177,-91.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>177 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>177,-91.5,177,-69.5</points>
<intersection>-91.5 1</intersection>
<intersection>-69.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>177,-69.5,184.5,-69.5</points>
<connection>
<GID>68</GID>
<name>N_in0</name></connection>
<intersection>177 6</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,4,89.5,12</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>4 2</intersection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,12,145.5,12</points>
<intersection>89.5 0</intersection>
<intersection>145.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85.5,4,89.5,4</points>
<intersection>85.5 4</intersection>
<intersection>89.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>145.5,-14,145.5,12</points>
<intersection>-14 11</intersection>
<intersection>12 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>85.5,4,85.5,7</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>4 2</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>145.5,-14,161,-14</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>145.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-4.5,89,2</points>
<intersection>-4.5 3</intersection>
<intersection>-1.5 1</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-1.5,89,-1.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,2,89.5,2</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>89,-4.5,116.5,-4.5</points>
<intersection>89 0</intersection>
<intersection>116.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>116.5,-40.5,116.5,-4.5</points>
<intersection>-40.5 5</intersection>
<intersection>-4.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>116.5,-40.5,160.5,-40.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>116.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-19,88,-12</points>
<intersection>-19 5</intersection>
<intersection>-16 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-16,88,-16</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88,-12,122,-12</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>88,-19,90.5,-19</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-24.5,88,-21</points>
<intersection>-24.5 1</intersection>
<intersection>-21 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-24.5,122,-24.5</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>88,-21,90.5,-21</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-41,88.5,-35</points>
<intersection>-41 3</intersection>
<intersection>-38 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-38,88.5,-38</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-35,121.5,-35</points>
<connection>
<GID>89</GID>
<name>IN_2</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>88.5,-41,91,-41</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-49,89,-43</points>
<intersection>-49 2</intersection>
<intersection>-45.5 1</intersection>
<intersection>-43 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-45.5,89,-45.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-49,121.5,-49</points>
<connection>
<GID>94</GID>
<name>IN_2</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>89,-43,91,-43</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-62.5,88.5,-61</points>
<intersection>-62.5 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-61,88.5,-61</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-62.5,121.5,-62.5</points>
<connection>
<GID>95</GID>
<name>IN_3</name></connection>
<intersection>88.5 0</intersection>
<intersection>91 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>91,-64,91,-62.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-62.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-69,88.5,-66</points>
<intersection>-69 1</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-69,88.5,-69</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-66,91,-66</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>88.5 0</intersection>
<intersection>91 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91,-82,91,-66</points>
<intersection>-82 4</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>91,-82,121,-82</points>
<connection>
<GID>96</GID>
<name>IN_3</name></connection>
<intersection>91 3</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-88.5,114.5,3</points>
<intersection>-88.5 1</intersection>
<intersection>-76 8</intersection>
<intersection>-56.5 7</intersection>
<intersection>-45 6</intersection>
<intersection>-31 5</intersection>
<intersection>-22.5 4</intersection>
<intersection>-10 3</intersection>
<intersection>3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-88.5,165.5,-88.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,3,114.5,3</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>114.5,-10,122,-10</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>114.5,-22.5,122,-22.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>114.5,-31,121.5,-31</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>114.5,-45,121.5,-45</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114.5,-56.5,121.5,-56.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>114.5,-76,121,-76</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-90.5,112.5,-20</points>
<intersection>-90.5 1</intersection>
<intersection>-78 6</intersection>
<intersection>-58.5 5</intersection>
<intersection>-47 4</intersection>
<intersection>-33 3</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-90.5,165.5,-90.5</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-20,112.5,-20</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>112.5,-33,121.5,-33</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>112.5,-47,121.5,-47</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>112.5,-58.5,121.5,-58.5</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>112.5,-78,121,-78</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-92.5,111,-42</points>
<intersection>-92.5 1</intersection>
<intersection>-80 4</intersection>
<intersection>-60.5 3</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-92.5,165.5,-92.5</points>
<connection>
<GID>67</GID>
<name>IN_2</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-42,111,-42</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>111,-60.5,121.5,-60.5</points>
<connection>
<GID>95</GID>
<name>IN_2</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-80,121,-80</points>
<connection>
<GID>96</GID>
<name>IN_2</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-94.5,109.5,-65</points>
<intersection>-94.5 1</intersection>
<intersection>-65 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-94.5,165.5,-94.5</points>
<connection>
<GID>67</GID>
<name>IN_3</name></connection>
<intersection>109.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-65,109.5,-65</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,-16,143.5,-11</points>
<intersection>-16 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143.5,-16,161,-16</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,-11,143.5,-11</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<intersection>143.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-38.5,132,-23.5</points>
<intersection>-38.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,-23.5,132,-23.5</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-38.5,160.5,-38.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>168,-17,184.5,-17</points>
<connection>
<GID>93</GID>
<name>N_in0</name></connection>
<connection>
<GID>65</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>167.5,-41.5,184.5,-41.5</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<connection>
<GID>92</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-33,144,-18</points>
<intersection>-33 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-18,161,-18</points>
<connection>
<GID>65</GID>
<name>IN_2</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-33,144,-33</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-47,132,-42.5</points>
<intersection>-47 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-42.5,160.5,-42.5</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-47,132,-47</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-59.5,147.5,-20</points>
<intersection>-59.5 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147.5,-20,161,-20</points>
<connection>
<GID>65</GID>
<name>IN_3</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-59.5,147.5,-59.5</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150.5,-79,150.5,-44.5</points>
<intersection>-79 2</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150.5,-44.5,160.5,-44.5</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>150.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,-79,150.5,-79</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>150.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,2.32143e-006,177.8,-92.7</PageViewport></page 2>
<page 3>
<PageViewport>0,2.32143e-006,177.8,-92.7</PageViewport></page 3>
<page 4>
<PageViewport>0,2.32143e-006,177.8,-92.7</PageViewport></page 4>
<page 5>
<PageViewport>0,2.32143e-006,177.8,-92.7</PageViewport></page 5>
<page 6>
<PageViewport>0,2.32143e-006,177.8,-92.7</PageViewport></page 6>
<page 7>
<PageViewport>0,2.32143e-006,177.8,-92.7</PageViewport></page 7>
<page 8>
<PageViewport>0,2.32143e-006,177.8,-92.7</PageViewport></page 8>
<page 9>
<PageViewport>0,2.32143e-006,177.8,-92.7</PageViewport></page 9></circuit>